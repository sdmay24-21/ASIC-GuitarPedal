/*
compression module

*/
module compression (
    input clk,
    input adc_clock,
    input [8:0] thres,
    input [8:0] slope,
    input [15:0] data_in
    output [15:0] data_out
    );


endmodule