/*
memory control module

*/
module memorycontroller (
    input clk,
    input adc_clock,
    input record,
    input loop,off_chip_mem,
    input [15:0] delay_reverve,
    input [15:0] gain,
    input [15:0] impulses
    output [15:0] impulse_output
    );


endmodule