/*
memory control module

*/
module memorycontroller (
    input clk,
    input adc_clock,
    input record,
    input loop,
    input off_chip_mem,
    input [15:0] delay_reverve,
    input [15:0] gain,
    input [15:0] impulses,
    input [15:0] data_in
    output [15:0] data_out
    );


endmodule